`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: William Shaddix
// 
// Create Date: 05/31/2020 07:05:05 PM
// Design Name: 
// Module Name: Top
// Project Name: RISC-V Processor
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// In this project I will be writing behavioral verilog with the 
// end goal of creating a fully functional 32 bit RISC-V Processor.
// 
//////////////////////////////////////////////////////////////////////////////////


module Top(

    );
endmodule